module Lab3_Decoder_5to32(o, s, en);

output reg [31:0] o;
input [4:0]s;
input en;

integer i;

always @(s or en)
begin
	if (en == 1'b1) begin
		case(s)
			5'b00000: o <= 32'b00000000000000000000000000000001;
			5'b00001: o <= 32'b00000000000000000000000000000010;
			5'b00010: o <= 32'b00000000000000000000000000000100;
			5'b00011: o <= 32'b00000000000000000000000000001000;
			5'b00100: o <= 32'b00000000000000000000000000010000;
			5'b00101: o <= 32'b00000000000000000000000000100000;
			5'b00110: o <= 32'b00000000000000000000000001000000;
			5'b00111: o <= 32'b00000000000000000000000010000000;
			5'b01000: o <= 32'b00000000000000000000000100000000;
			5'b01001: o <= 32'b00000000000000000000001000000000;
			5'b01010: o <= 32'b00000000000000000000010000000000;
			5'b01011: o <= 32'b00000000000000000000100000000000;
			5'b01100: o <= 32'b00000000000000000001000000000000;
			5'b01101: o <= 32'b00000000000000000010000000000000;
			5'b01110: o <= 32'b00000000000000000100000000000000;
			5'b01111: o <= 32'b00000000000000001000000000000000;
			5'b10000: o <= 32'b00000000000000010000000000000000;
			5'b10001: o <= 32'b00000000000000100000000000000000;
			5'b10010: o <= 32'b00000000000001000000000000000000;
			5'b10011: o <= 32'b00000000000010000000000000000000;
			5'b10100: o <= 32'b00000000000100000000000000000000;
			5'b10101: o <= 32'b00000000001000000000000000000000;
			5'b10110: o <= 32'b00000000010000000000000000000000;
			5'b10111: o <= 32'b00000000100000000000000000000000;
			5'b11000: o <= 32'b00000001000000000000000000000000;
			5'b11001: o <= 32'b00000010000000000000000000000000;
			5'b11010: o <= 32'b00000100000000000000000000000000;
			5'b11011: o <= 32'b00001000000000000000000000000000;
			5'b11100: o <= 32'b00010000000000000000000000000000;
			5'b11101: o <= 32'b00100000000000000000000000000000;
			5'b11110: o <= 32'b01000000000000000000000000000000;
			5'b11111: o <= 32'b10000000000000000000000000000000;
			default:  o <= 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
			
		endcase
	end 
	
	if(en==0) begin
			o <= 32'b00000000000000000000000000000000;
	end
	
end
	
endmodule
